//--------------------------------------------------------------------------------
// (c) 2022 OA
//
// Module Description: Timing parameters for Hamming Encoder SimEnv.
//
// $Author: nebu $
// $LastChangedDate: 2022-06-26 18:45:18 +0530 (Sun, 26 Jun 2022) $
// $Rev: 21 $
//--------------------------------------------------------------------------------

parameter t_ck = 1000;
parameter t_s  = 80;
parameter t_h  = 50;
parameter t_cq = 90;

parameter design_latency = 6;
parameter duty_cycle     = 0.5;
